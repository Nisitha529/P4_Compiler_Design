method _routing_add_entry=ingress._routing_add_entry;
