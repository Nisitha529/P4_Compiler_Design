method _routing_add_entry = prog._routing_add_entry;
