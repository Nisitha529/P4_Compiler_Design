`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
IEQCf58ZmsaoE/XJ5HZIMNJ+3454/Ba27Om2IelboUGdhL66OUbScUzJkbz5Zs/JL2tOpTWRbPFX
x/xwukPCnDOVpNz05Uy58BGhRahqx1yGA9JopzQclS7ftnTx/SeNxydbpys6UDdpbe69GkU3VQyE
pApfycr8HlX4+/b2omFUuTPmzTNon2gH3999P7MOquobtQvp8hiF8dj0hL1FdBqDcI+KBzpQKtFv
GELJE4NRMYpxb0x3wfZZR2KCotwf0pv7esbY7SGpDk8Uo2vLL5h50ANfiJ4xEn0oYEzj83EZer/4
yb/Hj3sAu0STs3mTAnbaaFp+Vwst5xsMEoRY6g==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
kHKyfyH5gm4S3mDmrU4ZXZYawXcgDmuEq5v42E8bbYR1L/HrCQuoOup6Qml0T5xV1JMR1hmqGyT5
krEo65BfLPrmoY/7gqsL5eJfbQ/D1HuHt/strEuC1XYSPGdiBDsH37xy9KG67cNUv42Z0oEt1Gjq
3TK+czPti1pq+nV4FpcnlzeOBeUNCi67f/IAOVetrH5R4uKZ8l2a4EKsBppK13q3UDMoj9kAfAET
X+B4g6s9PKz2WCsdJiwfl2vhQCf/S+D3h11zy8r3XA2dtkifZE0yxE9x3EkHYXQpICBfaLYJwACt
1VK3dYOSD0qPKYuvF2/wSUkYHvgvhmKkeOjKVAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
koZn71oMk1jLoNh4PGMpBtc6aiYMflCZQVIlHMqI8mLfoY14W18AzgqRHPN8W1ujL4plvG5+XB9N
Gs/Ce2v4cg==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NWC56T1dCfCj8Enf4MSXVtWQv2Dv/f+QwqtUH4yPihXTSMgPVOhdwAkJONQ77Hx7d+FuMAapZ+OX
Ejzw4Ml7B1OMUklFaHL1AApeha6wJKbkNvQNc56HXl9ZhOgote0wun+EpWimwSIiyPDjjGmd89G9
fspSxl7SDAm1nsEQWBWiYlX5bj9fNIcNmvWBSqLCEqwdvt+0cQG5oCiTy3MEUJUHbzPgz1fq0RWI
hH3h8yqQOLnagqwF9PeasQNfJ+7DT915NIPsDWgwF6+/AxOZYgyZcRO6rZ8Wiwdj1Re11hl9L+We
ETkpg8gMYAuogZ9dHimPEmyypbXQw0L+/8QClg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
G4Hmmazlby1LazqStVvU2S9kqjl2Tg0BautKwetSSyL92N/SU6sn4wqWJVs69OAay264FBWFrvoM
Z4IJIMLfcZLKphcH8qWRG1AdAOkeIfTyj1SUgzDWbTEMYzqgE35F2+FSv4kcOnZSZaoj+hGjX2fv
evSZuZWwGqOWJuVL7Szb2QssnrsG/40gBUz6NnjHh0eTvNsow4JjHp1cERd68CcC9ncjPCAr7QLX
NzLNRpRYqujbRXHb2uA9nFWyXkpUDEu8Kwb0b1xSM+3rSTUSKEjvcy1Bb7zeYnGPZ/VzUPWid2vK
lOKm46X6cnFz20WzW8bvsrsuN4dDe+3swwuAlA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Aw+kFEVQYT4VfsPpA6vLlqN2MDy5L1QNjKJjlGGzTzLrpVSuOWoPgxLTr4z1TDiWWDfbZNgjYNtN
8Aurd4w7Wb5Q0FKv7lAfG0BSfCFWmsN6UM7TaFv1w3x/MMoCMh23Zma+9FF7MsVh4hPfV/9t9wEa
d2N/DWIKw3A8yF5Q17A=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
q/pPD0hSm6ZWKasCdhOc1oBa/nVm30KWZwDp6wyN44EOS7JMunJL+zEQj9SEklRX6mv000R/ZXnK
CJttkm+CmOfLemxWO0W0XdaX3tdjjbln1hWT5jOx2iTmFHHW44FYtMrWQDndViF3PPU5ziLHNxpP
rR1zF0w3pXjx5Bb3p59zeUbLJTmGZlD7KD/Ou3h0GpCbRDi1pVNs/MQpx6drBnUKTbbo5HeXz7uT
M0BaNEvCopLr2ADmDZhiEjrQVTx3cFSjj224H3VsTSMYTu+7hP4cEIYOx2Xtcs1sKZDJWmZV22D1
VomiNGlEDZpZHTQKXN0uLQCrzg3lxl1Uk3/bVA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mUVe3fX9Xz/bkGuDwOG1BA4RFiG10brAalOIgRvvNy6lqBGM5mDRKk9TfeKQyyafH/mfsULMVyaJ
OFeE3yGz9TzN9jHqM6eX0iurKzQf1QJ3wi2RDEeFWMUX1Lt+in95QpfNpZgitk8/1SMpyNCcWGNj
PiBDR8g+Ke8e0rsSrCt8qsAJO17iHkwb7zdBRqomA7ffAxIkiIbhzVDU1Roi7uq5Z/MYII4G1qeK
qtJAn/3SMp+yzAuj+qElIlsybGfSSsOnHYXXI3I0T8v23VGVoXQZjHAwoktJ7NR/j+A3V2lOCBow
lqz1yk77QdK4QsupMb3uDhgeRX2OXLn7WTJZKw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
MNDl1pvX/zg5YDreYaFBCnsJ/zFyCGv83eF2JC5pkZ7VU1ogyXq3ZXM8xV3CoDTsZ+wZURAhdxpt
xlTvn3wv3Zs49NTkxpbfK1On+D1+p/gadT8jS3vUQIOVCWOkN4DRcI4ZAdXrPWpQ0wNIospsy+ej
3Bi7ARKOlv6nqA3Gxvw=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
neoWAkpfwaUc0uBgiVBbK1JtH1BLeEl38NG/YcAmhZYkQJ76VcIQqEZ9xWr/zm2DbHCZKLlpGilV
oaAdX5zT2L7ksm4YWnXroiXOjK7Sdi6v8LoKAjovogAzY0GJkE3goR5PU94RNF55oiSV7+vdU6uP
SK1igXjeRqfrQkpKLhLyJBe8cn6bm3Dv4/iNcEy8TD8c8htYHPMqpScwKVzvQ/bCjiKYGA65vWW/
7C2ByDMksxp8O2Ada9lyu8jkxZ/b7JnyClmAGgR+v0IVgMCnqXLGFULhY6TzXB7+YQkakAjpv/nA
q7W067vN84P/8Cjh5u77kmsWssIZJ8mkBNA6NQ==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20560)
`pragma protect data_block
pBn1VM7/50namOCcJ98bYWTMZKcVizuOow+vYazDFwfIcukpQPZ4JLKtDc6JMkRxejtzfQ2i4mvU
NVK8BAkNhylx+ai4gGnOee3KaJH0FaX1Gz3YWaD1Quw24WxVCg+yYB9kvP9zZgoEfMv75YHQxMUg
BgjguH/Q5+mNrlvg2P8oO7JLe3uUg6EDa2F7rL6QCHvfy0P2ieXjT1WZWY2bMbR/VXat7ugmBRE8
FUgP8sJ2m5+VzzsYmfV7swHZfhrDLvyaLLjuiTbyF7kDJLt9Wu4I8H4KfaH4JKBKdpwRTY+/Umfy
Kanjs2quMaTBvMBf5oMWqfFbbHCSrdtNimt+G2JetiOxwT2+6KrKab50GfS2KfVtzKOWBgS9nOex
oaq/flwNH7NvGVgvFLHoRL57Rve990VEDG//D60WsBe2Lp/3Frt9jLWI/zxjiDQh3ARxGXsrl2Uv
pn90+2756Qjg8qer8GBgWMIf6BLNxm9zAHFL+xehJPvHCAvN87P/WU2XsNAd596cRSofD/AHBhMK
S7e+cNUzpgFcNibIVLJfq+S4RBQO9HRhfJrq71/ROo/HnkHSIzxhp9xwDS6jy+vXY+DDQAJ2xHaP
PJ+niH2pNDqaUcuifuWWS2M5qxQ46H4fJQgV4X8/UWc+aNeaClwqc9GIZAgfi8Ofvb4xtlucjdYX
gPpUUN2/3buchaVV+oFKtm5XnIaQ+wl8054jdY3loAD1tzmyymbgkdfAP7aoC/WThkNhU4O/SlKG
zQONV5ac3q9A4L2z6PFZY9/x+BiJX0TqUdLk0eSEb7tljg45fL2tY0h/m4gi6l07kcixGeRuSIVe
ydHDvR7sKb7qlK9Q3Z1j7eO8p8CbIATaTCPW7BKHy9kgDXW0ACOSeeH/wqiyaDsDQjQz9JhEFGKD
Yg/oRlC9s+JdcFXNikScyGZr6JG5dBfvJqfgnws0IJ30XkrSZU7OC8bCA1/ozq+g0JJZCC8jidWh
bk0dJlSp41ZDqvvtIgahZBz4qhDd6LNLLI8qt/bo9877izGfTqcdn+YhT18ovUhQ+NMTH6aUO8qk
+V4dTPKq5upnDpH5Y6AW6nD138gg1uEAbEfb4AstFWE2qRNuD99sbIRseZD1+6pPGNAwN/cf/BsU
/POcTm+RCmhrCosRlHRqURt5Zj/+GEtSHFXqOQEfz+KBSFGBCACqNY2CGse03qBwrlYk83MGkbOF
3Lc6nd2ZvxKxSC0KKgmxn6mzinedxmkXHm9Drpj9rCkLlO0Arw0mIL3ScpVeCx19ELJg1aK7ovbK
CSExYFTUM7q6wfA9Z7zy9vDwlU8Rc4H8hz/QDAmKW9gdNHufbP9+BEjFwf3AaBpbGoFM1EO0+jqv
/STnnfrl23PvZzD86DnONRD1CbK7x4EqqVkHMRpRQcKnmYrs6dVGJR+oJ9N0VR3R0dPw3XgqKzQa
akCTFRihehs99RVJzT4FZkV5Mv78NrYEFg2FW/6L46pqJFSsdziUmtQcnFQ2ifZYDXrjVkCTKXwZ
yLUqOG5KAGd4vCQGUFhMPwvP+IUBvezyROMu2U7bAIU6UHlROapHn3wiqvrWEtErNwLT7q3Fuyzi
wp49efRI40lpuLhPXZdwGDkIOuLnE2O0bvHSwVt7lC/9I+KIO1JtzmZCdJsjHJWynW5XqDekXuW/
RKJP43X7d4LBmbpRk1Y2LQR7vuPo+9vWpfTame0L75KEgTzvl3e6yN5WBd3UPPBa4VFx8zvCiNS5
N9OoQBaClQbh/UcZxqG21xItYVvNJ0MC/53MUzAZ9eXlD7eDt+M8fxIGZhWJnxZOW6tA9Uiu/sJv
gEREUXYwy1m0+eZm5gh1XwtODhgswAgN5fgpgzLkRHm0i/froi+YJm8dRvzkcI5RnCyaA9PA+ZL2
IbAtqm9uuTC6A95MsWfSOJOsN/NiNdKesDK6p8cEsrIKD21Pri+CrZzPlE1HeNguaJv9Omk11H8s
Udve+TvTJBIMOgrkwm2dnaV1MECph9ouojaFfKcs4EjY98Mf4wHN5VmsD5+ezy2gID4UNywrpnsX
qLcu5xsPYiKF3icL1GiTR47ISPv9Tr/ym78vLzfJossj5n43LEiocY1QfUxJwQQh4UBxhat27EXf
LwpIO9gdXJMOjeN2ji43PlvqBJIUKYEIfwP/qoQ5NGv/2i6SSK2yFVas5DHaloiRn7T7M6iRHcLx
fLEBrllge4KtWkmroi/v4XQprjAMp5i7Z4hfcr3T7nUXf41jH+K57RR9hwr62L06qVclDao1ePqm
Rta67J8qk4obsFDQf7ZiVtQPJTw37p52Qsg+dWSbjQaTEezR2jrHKgxcjsubc83Jp1uWMydr0K5F
93nQHg48bn44vGMQCwHUyE3ijy36KuPVcLOEI8y6Zs8c4lvNU18SEJCFetc9xyJSZKlqD9S+4x4e
m+/SKata/dT37FajBIPi2+PmtESBgrRAX71Ytm60QFyCYnVnF0TgR/4Y4lKIc1rgT++cZmx9edep
Vupbll/xk34SrVmS8MtWhDFWTQVB2dv26P8CxfWlaFIJuEzwBGjDAHKEHKT133PuG8Ztjolm0ZkQ
TGPW5iSm/ffbUPt4BoRgu2lFqyapDLsIAa6YgH3pp9CpJ+BjygGy+ILKWISDLcqy3O9CO9pSfZYD
DTThn96fI7w9bMrDd0JQfiT6wbHxbjkF79LlpAMOZDkoO4Lj5LQR5pZAalTle9QezO7ukwhi2C3j
LQY3UFdrJgwhdpFXENTpZUj9Z/M+LQ8fQTlFEWmBfhXXjyR8qpazIU1xlwl1ldkbsJpiQ5NdwmnI
Zt23jaQ2zrwhYC26Y36PO+rFhncTXS7kqBETxMKm2I9TWUhhb1v98PX0NwqvwolGTi39KYDi/Lus
qiV714F8r8NIqbB4C+rE2kN1wQ+3Vx9dkymT7A7I0wBGOEbAfKdLfkYfL82paZbTmXcScQmZCqa/
ESKPACtr3aHXmF7tgAkBZb9OGvyZ2qoXuPSNKZt9vV5fNse8+QWrfEmMXv+xNQiJodZdp9duLTeq
1fuAJnYg2eP2tEeI0Ck9ALQ/R2XdrwSz1/24TXDSRpHZyZy+lDn2AtD1JRbJ3M0Ca6fNIxGrcXY/
58sq13/QeHm1JLB/TnWRqr1yTANf1cCVPcnWln4vJTe2oe0if8KTqZmE5vdD0cAjH6e+9N/NGDes
l2JRxtcZ++Ja7lC7iok/AtQ3uUvKYDIjvSUs45yEpOT7/rc4wts8GMsLOPqq6ANzH5QAxgYIgqRH
U51coQvJwB6uTvhQaD2jgh70PQg1ns2IP9/CxNFOMeiyp2SFh9Je1F5Ezdu0KErPjqqp1N8V3/Kh
2tbmp40p9YtSHUc91RJ8dvnvHaV2VhiMvwPEf9kUN17LxDhjL2GxEo+RDgJPClo4H71MBMDO14J8
WLLuM2SsTCpBIWrgTVNsUrTNBgZ3neU2bL0+s6VoVi5nVSjzwyLVyy/YtAgIQ7dsZITczbH97fhR
Qrn1WK6dxPxEiRNUorsQfZVHUi8qnjFL14LM4zIQBhm9+IAkFZC1DsBofEMYvMPhq77Gs1ojAhbF
vmRzAbUH1mqnV9xVM7zFqkE0vDL9U34bepcGOaKEfbChWJTN11EbFvpdjxw6So9zeoO7uHfj1H2m
+iC/GQH+GIxmjtnrq7S/rEk19D6Hope4DvOEC9W0/Du3iY1nfSHrlG2/J6kqopM2DXUP/y2NOfjp
T//xtGJoieBm29l7Lwm9DQ16TUVc5rsyIV5TzYsyYrHVtcYb1eQJgLUt7GYa0JpVmI0KjxZovKjY
1jCPBEm7r++0h/XxoDfsZg9W/Bj1I+4+tWXjti90eb5uPySjP6SvmqU+ByQdAFl6zeJaoyBxO52q
zNEF+KI6jt2B4j/o8hXFPwOspJTkVP2SqbmBD+VGK7NzSm9b5jVbBd0VA11hOkEHXDGq96AhrBWY
WgFADlMXIdwNWNwx7osBR40fJDPPy46R/xgrZs4d+TwfR7DQmP51yKC5W2bDzvpwdIqGcuNmP4Z+
MvYhvVb6lIcEWMzM4qS+428+g5oqsbr8wGHMMTKkADmt+Xy81Bqafx6GaDTiyyVqifc+6UBOu7zr
dcyQdg6YEIOZTqP5Pt5meTcAFuH504lwbLdYt9/cWXObnkv06XqaOPwDzf/wtJ3WIxlY8t3h5Ym3
/ZmtvLgYXMrrncvGLqWsPSjMwWq9PhTE8qhx8M9qzNuSJeaL6t+T1I4V+kZS4KVItFZztI8UMvFR
sNJVIhp/3yNZCfEiC8dtFgSsLu4ZEBZngzzun2EDsSTwR5LXg1Lm+UfbPCdAGv9/2POcPUqlod2J
pIL/GWDa2QqZM8HjvahmjOFmweUac6fy7hErOGbCQcWXJ1Vz6xYyZj0Tgx2xVuVfh/rpdyl0cZbX
CXKYW6daPFSB9Hu3vFJs1yylASG0MNqu8z+2IY+1oDYm7PryXRzhjtyKkKdl8WhO+ndGUVTLFPN2
pHfQom5YEHu19MxDG5IqpMZrdL/J5/B6lsHo0s4ctLmVkP75dIKPv32NqA5Aw0MshEi4/sl/Pox3
DkhRWDUrG2Ta8X64fIS4l9bYI5cXo45RN2Vjh+kEZ/Xbe471n0AjrV+8GAtGInw3lj9bYp3kszYX
6VYecFbbqAQxfasffS38NUq5qlekQpznhrOqiwc+CQ/v5xcb1O6PP3eGD49iIJrQ5T+Er8aWy0+K
9Xzk0oAbY/OzwvNnhZwNZEXuAXn1hykvbtyHCm9jft8XAC3zISLTN1WOJDSd1f1/DIWe3O2hEnZS
UPXAjfQTK6E5wavduJvi2IjA3L9YsAHbDfSKXWdfxf/R39YdbZFbVryy7G4P42vz2KRU/Ug9cDCO
7j3bRd7dYYljxMrAh2oY1/kHVOC0fdylzToHnJMyTdzrCXkVcgSqxpbkY/DzeH3i6waxoan2ZNiT
2sWZ7M4uiUbVGPBD2eD/9MQ7AYe5qb+1535/IvR/LelcIPC75ucoxOnG8Tna2MLFuKB9ZeXDOxFy
Qgd1HlOYGTCJde1kwxNJZKpn82Lq4JVyOSaRz3TqHH7noiAEf2C4A88KSEDbfH3GGwYsT9UOI1sx
HzhRJQSK1q7YDUMXTF1v1ZCk0lgP+Ne8Bgw9/W7XIAnR5oVTfdeQX646HvGPAiaaT5njsMYY/E0n
6l5roWk41y9a8W6FRlmsm0xiG5t6TXTBCYBvMWOu3627vFWHItYZksRkrhX6RGqy5LY20VR8NIat
8Kn0qFl3tmmLeTub3kEDUZePjeyYK7fhGD+U6Rfo6jG0gzwEXb5I+tcek70NGhdKYiU5PIx8dA4j
KY4mpd1v7ASb7oy+bFvAwkPIa/iWR5DZMVALvfWqQxzQ79PDn6rn8CeTFl6ljNqVaY5S4ur8xPD/
sXU47jof43041joNK7fyK5Gv7j/AxirNNERHTsa+6BgEKk9zjGw4lhFoRUsCxwSieo3hWF75yu4+
Gp5wHkJveAXMjx01fmKgoAIhr5QwxHhlQUzHFHY6WfHSu2ZBJqsvA081D5agYcKS1tsQdeUfj+5C
EeJ1nMeQApBcCd/GW7raEXpL/WnSEuG0jx3YdN9Q/2/VQksaJ6PwPIe9ZHzWVLT6j8LgHi8Qp9oH
NzqGNO2ylBrWAKGdovEEMbwo18li4pj9iiexthkxn5JJlv/UmaIK7NNGqGH4n0HuQ2ohkbbAoZ5+
MkLbr1IjHoaN4r4ECu2KjJvB29uSYm4MXC6ytw34aPzjqwut4sg7eLbb3WCFRywg+q32/ydNUJc6
le8icgGGNEVSgYJ3JTzVNuiKp2jafX6fUrBEvLwCVHvcF7/mZM5V1zuDjTgKzGQuavCeDmjpsAcN
8ew88APMg/qU+Qqv6GO4rvakdnX0jLsq9XscTjrbLfipcNdDZZHH0lIDRFmsJZlBSjS4On3MWj4V
kFH13PPG0RXjPMPgGMAS9R7EXCtu52ZdoW/L7qeo7010XM+ql6/tiRwahuuWcLUsLimwsENMua+5
xvEYPIRVBmz+0xRSZJth17SELdLEg6yH5/yqgsjt5LYX59eBXRWoNQDzVBPxrXSbbbhFppJA0tQ7
BY6ccF24xUVZ3RLDRl8yA3l0rZp1Z3GuLaMcCqLrY9wdlWO24Ypre3SqNDCp57fPG4//kd3K4PYr
yBL3DSgWAf1QQw+osxOYv2ywTumFJcJRxXfjKjP8dsnyvfNBA7dYJ7tYuKSiBRsnkBql2763ZwUv
AqD5LtQs7pekEcQmINc5RrKZ9OsYW1F44GxgiO/3V0WwnxF0pyIC4WKtC6inKv0S45/YEV64sJZm
Bjs7Uxnwlol1B0Rfv1j6zh/WzYxXYPo1JvDsISQA+k54t44Kt5dFxGhDvvaCTqSOaQB7AqC8tVgZ
jn9Z/gSRnB0lqwcMp6cnKfUhD59VHSYPNj1+QnOjHkYEnmFwMUznCC8o6A2hYgL4/wo8NDKoTseF
MIJlIoyTk/ozY2nDZuBTNHLXEOHl7HZJyReMCeCVeyTChEFkV57miyQNHPqeOZ6JA2D2h5SQaE3j
vzXr6oAnB3Wi4Z0xK0WZRB/uFInpcQRqLC5lLc5PlR2G09uefBG+Mhn8lpkMbwT/yjCnqnLOB6pC
AMxQMKg8wnKcgNnue+6txuGZMB4hJBjYelIMdDN8RNaDkhd0IZO4rYJL847BrfnSW7171FAzOcZT
XdrzFm/JoZgZd4F+6u47oWC8NCykGIPRO1mak8PXvpv25iOkW1AqrT3JzczkxZ7kd95U/uK6yw3o
A+7/8/p9n+oWjhOlJOiHARc/RzvBM0qptmiuT09ghfFpMh2mC5VIWcC3OWRavoDaAzwuQmiyxDjw
c0xk4juw0fqqvCwRyHMlZ8mATF8bumZsZ+9fJzTSpjJNL7pxQEPg+Q268wqj4hc/6q6WGyPxREVl
omaV+8VXh1W33fWB7ZfW7pUhsBVeJzUpUPlhMklRixPh40ScV+kwtZGf8Slnk7tLv95iAUWV3F8y
lZLJ96Y7cXiNuoLYPphKfJr3sSK7RhedzubdK3eQ6Fa6VnqS7eqzSUoHdUMTGjObWoOoymN/vTIE
OTsQ6YzrMRZxUXOz6tieIGOepGZgGB4qUFqButramPGJP3jegcCjdbeQAVDYM/oK8iw8spOQW/Au
/tT0IK32fj+SQFlnawfGYHq1xRbhD2jR8cO/UPm7UVIdBRr4FRCNsCwWbBugG4sRSGF8xRO1s8xt
ibppC+Vl2yeQwfpx8obPY4Tw4beHs/GgGEXKxKstuFocwFyYy0m5cBSfvbNsbNFKqvw6m2l+mjpL
Kxd+FFdp64h+htPA7qNuJ61n6sSUYYpQhXcP8jMAz9H8ZIs18AekhS5TSgR3yHvwkN6sa8FWihGY
Z8ywCIzGjrRvpRTJPTRovnD26dj5/lWKPVxVCyff58Ge4mUrSeN/SN9DVSCYJuz6DKzFJO7Q1ciu
pN/gtBsqi8sW6SYMkhzKSVKLLJyqdP7p3Ig6ISeNI9D9aLxNUhesGQUvaz+niXdecLUN9KEkPJp6
wntgu5ywftCFEJt/0TsNHMu4pXK8YRPcTm+4GKfaFbHNE6C2qfAxzF+nPaQchB59/DfzY14ChAyT
s8zy1r8kZRw85EMZs4y3GbgwyJtgbuRQlwdURjBpxdGv5k0j5m69I+RP5y9SAV3DVO3meV4U1Pzf
izETp6XpinKZdw84dSz4cBULqz8r7TKj37CaL2jP3Doe3pfYfpBXR0qCsWEKiBWI25hVQA6DOR2b
mOIUpt4qrQuhNfgYNOUsH2CFcNb+nAW8uuwZgxMYQ1F/m5cm/+lUsdNUfj+tAAoSnc+Roe6Vc4Mo
/asl5xRzF+zOdu3ZyK4+JcN00ylMJyw6gL6SUTS3oVUCxxjIGyNeq8vOyLUWHFPkLQcmzhnnJWU5
K9z4XQ2ipRS4UcAPo+vTQwTvCC/UU3VY+Bxgqo55uQkSR4dLzHY/V1ylLHUWAkDtmHJFkAsLg7dA
BDKS2/fltDepwtOI/Np8dqlsYSHXku2k3aE8lUCRFHXYO0Mx2GHhAUvDwQL2A0yxig+6gHGyhQiv
VvDusUhpploBm+CV+h1+1qhn/mx83SwNSacPFNLuz/JKuYAYWr16EWGuE+WM/KibLwn32/3w7iXw
nI6+/uaDFdYWsBs9ib+s8H/Rhz7jYvzJ20ggBx2iaf3hm5419+6EfTc43B9hNdIC4RB30+3ZC935
fNiZwZTidD1zU0EwSXyTCdCOcyYiNxhhHAxtDJrtU+zk7O+HsAJX1mjwipqqhaCfQFsqfecRL2tz
0cdJrXcnJ94FsgRGuzWmEsgK8+GXhIpewhPlwkXH4q46Wb8PQ0q9A42oDhwKekGYl2XocRQVwuiY
0wNnzkLryVEQ2u9qpSIt6rS6Jn/INu+MSy9n/B2A9lqUYCHHfZYQ6UORDPvf/MRb8pYU6TG6ORqo
UvFQf5f0mmk3XkUuTf4UWshPZWLQGBWBcN1snyWbZbxRh2HLxnM4yO2i1tYiT5xUTX4wcOIVc8F9
KvmqGBM2Giaf1Iq3953VU0sBmXuFpXP+la2UE3KL8DeDvKzZjZizeiTkvw2Gnn8tk1483mEjRcgA
iXRFmip9JXVMSBWj5VJ6KBGZByE+JAKSDIHZhPxbVKeW/VwDE9why2dUoT5YSU1f6Bqh/jI82Eu3
OgoLtthB2dyN0nGhXoyYZNHaBKtC4QanckJzu9JufRvZSJv4LPjx3zx0DfJnUJh22Owv6xHBw5xX
7BiFxEpm0P6kfD5FpJsxYMGMnuyaZ06pLD4BXFlOC8QFWtvYNslyecSAHL0wvPG/GeV7C7QcCx27
eVQU5Qe3/NyaA/2pQlvC+9XXLkV3WjFQLrO3EcBA3Z2eEwU18Ee3u273O8dj3BpzpvkoZD9/tGbj
Gv2++J0nIx40ajyYh4WaoZzsrOndddJtXB2XsMTwd1ixAcBA+TYtIJKgE5Dr1yR1G3jMzV9mqXJJ
LH3h/KLf4nJ8f9kw+TuFzCKAKMMKA4h7WVoxb2k2ApEQNPoSMBkI5xuocVMSqi2FMs1IEHteqwKD
Oh45RCp3znOiy+wr/aZlZcKG39+d6ld71Hv/+ncdn4urNt5Y90nuCUeAsUyfzGTGArUiWK9i0Fdu
iKEbXkMflKLrTjLOOphojcfd1wmb4iXRsdtwhy9kowUbIpwqAgxOvyLV4NupwqAL4zZY5IdrVZM0
1+97xgbxzA644DCdRCcgnmIooVyN7zRsTnbsJ0B+s687M7dXrfPhKdlnx7k4APf6i+iGKRYJCMSy
kFMyXAJER0cvmGTMZNKI2cs61ZVnh2r18VN8IeyHnwgBU6nJa8zCbZrMSQBjaoORzRu8V4q+7jEP
Ojg1j/2yXEUKDXUwMp+cEHbqVJoZthDzWb5w7ZHp8jfvQDPN7eME6gUOg0hrJLZNeUvWfvN1Okei
9sLTSzp4xwVR8G31cc87p/S8jUOPxsVONlymHl6fWT5+ev+YUkaoFmWIhQ4wgv+Rxo9YUuH0maNM
GHPTReFHg6CivbaOzKRT0JkQa1fDLEmt1FxR56xy2bx0RBci6ztDqrQGi7n6OvCX3qN44r8zBy8M
pbPgXO5il6v4gXTHKpUEJpBbrK+haIASR9hzybWdlMjxHpZyexTGH6LU6Q4eXn3NyvffKJus3GLb
/fGbtp2TWsBH+x0QWT8rLJaOk4TNSR5WYNs1ng4V8om1zqShijqtrcokJjWhU1Ph/JSFusU1Puzo
PZxsyaTF86cx1xYg7L15ND10VtLHhciwnhHLUTPU30qnRWbtaMsPBPO0m25Tn5izkYLvdzDcnbwW
GwMW+oqtFlF+ygnFSO4QxKNzreArVjr6DiC5EknFdYh8xb0OW2GLR2cxeEqdvObxfKz/ju/eSm6h
0Yo6hRfOLmvzLUV8gnknb/X05KRuE3UIr9QVFhpd8o4C7Ag0m9bXzkP78QHkuIXkDaKsHzhccseO
GlwpxPXOgtKP1wevnOkRoB87yV/8MLIaAdung4Rnw1+qxe59So+teSSZYPoBnvke4UE9L7/3nGnZ
dprhJPV/VKvCMtZ7ImEXxh3ilNQPc9wZiGkjYtvb6PWEdK8GB5Kr7Z01IL+SIhxHWpp2oS0p3J6W
ZwXFJXk6473LaCfBwqUu6ZKALaTZGnTJ1HMa7BPkAdUh+oH2bcPopr9dw9uvGDuFfgdHEEt7Ti//
tmIfrjTmiV9N1sdNUrlmm0+fPSWbw8Hlc5eJtWLVl3vWdB9E4GTMrmZyIkcQvZtmUhLz1KRl0igo
0Ir41ezQ+dkc5nZYjxPx0/QVRiqMjPBElMS6j596BmHI2iTnZEzLUg0JAzCj8nkOxW1uQiF7Jomi
MSmbRc3cIePNnTJoz68gC7fCi/evqsbFJCsL+88b+5FXcJBRgBqfgjXCJMWXX+vo3DFnOSFcTNwi
jN7UGsmBGa1ycPRQxKsMoZSoqcB7+5L5xAvVJRn6ZBNdJwGJOa6G9KbvLwOIxdrbS4pzFx1TYfIt
myaDRwgLhk2IxS0+orZaBn+zJUeI6w4Zw+6jkwXpGfgdxynOaYpu5tk8hblrW5xpE7kgCBfvbF/2
awzMMyvRK3qboUG32SwIjqwoBgsWMxrWrcvdAkLK2GvEysMSEVQWqE6rweVCR4Qpsylu5InnNlcm
ah97gBl600BOSG54uCsFfUHS0RRGiyMXznTXJb6KQ8artI1Ko1dVDUP7VV9NhWmvzv8UK0g2NCdx
BFFsTbAr+ZWWvkObPQxJKySLgjpcSkZPVYa07UA/ofxRhEybmMGegkWoXgU6bTgthk96WEnMPFpV
rNbxJD/SqMLGgO1suK32zzzlNrn3gzv9eF1Lm/QdMx0qsZc0/qpPHjTNd4frVYRrllEINIOrvBsG
OgJdZvUt3BG+W9SFtRHCyNxrbIj1JkSFSPwGXKsq5LmxwGB4cRzupJnpdyBkfAlAhdRXOMjAelxU
isNwTo1vJW897g5In4Rur8vIaYCKxyYc2YzRJcw07yeFLqnKvieVTMN/vteXjXVQq0i/mBEqVI9m
69LyaAUSu79VzOXh9oadUIemJ1abKkM0tSZr64ZrkA7ZFbu0+dcSCpM1jdr3c8OcIFFFS5IXmC2N
hUZ8HGrlp+gdD+nF6c6y5gxG6Obf9FFxCcVlyb3ouX+0oovQEzVWPw6TPVkSIWBHVJIwr4+bveuh
ep1OERNWDlCKXRxiHVgyW5ZEHeXSm2mTmJ3Pjh0++APW80mfXLDcruT29F+TuiYBa6cqykh5LN38
nubw3Ljl4fltXT9t0rIN4QVl55DKkowceINn7xZGUPPPa7gRDoOMME40jRMcPlGRXUpAq2dVgiBo
O1v40gx7MOIO06LMrAEiL1bBKbUkBeyYhOeYxFoQfLmfAL9USe1KHeCaJzpTiplp8pW7676iErdP
XjEhc40IVK6xK/nyxq4fARf+X7EfMxtUBmwCgGfB6ZsLpEbMqabpHBysQ4b+rHpz/FPzLgbE67+X
DBxg3+ZGw/jC0gog80/kGPP+CV1v6IYqJwk6TykScsrmBrVKjRFqDp5tRP8ZhmmnjzOFfad5DhHq
4IlBu/f82r1qmqhTt6islLG+MKLAcEKuQgo0CzGsL/Agbdh7wmkfFXyAW62mqTcy8v+wI5PsgCm8
VYjBk2SizOfmnG0PKmac6Ij9bUJqiATZHDNL01GFWB6uQo53g4SdydTFHnikUu52mvx7k5ADWHZ6
wuIpEv87M/822lqzyyeGqPgS/IyuQKZfIykl7zIzHVsh27wsiZOhrppdZkpdHIQ06uXJ8JUq2phJ
bS7XoYQBQTfbTNDS3H7XYoIU4wPxS01MTRk6RYLHpbBclIbPAenjG5Il0nHR0lGRK/+XMf6QteG5
893ZqHUddHCToFz1syr+vVG5I3+mS18BrFlGUb369OVo7D0vRm1pB9UJfojkZ8ZTY8H75FS1p+gO
P+b76UL6tGY78A0OwsLQQX+0782FDmMK9oQzLImKkRRsq3LBLalnn8xoHxaXKLysbiTUU2Lj3gWH
5MqMHEDbKnWZ+biZWPr281XyZheVfxuepPheVXIOUKHyZDRy81ux8rg4rgQ+DUAKqsCvHs9E/Tjn
rS3tRYaVuFEHrHI5MYmsv47+tYfLHg7TPLJSHybYgWwTyNxihVP90bFHNKcdYR9Wg8XbXItX8Jyr
TTbViLBVqWDjso9GnTKk3t6Vnxhyahl2wr4LU6SnAx+2W0LRCWKb3O4IOsB267bIlYATYHZGwrSd
+38Uj2hyzkxePlLekLC8cZbPha7fMSCRs8IKZtf/kgCvoH39XBRTfrlZvhP2HttxgeCdoeP5qwjQ
OlMc00jhv7BhXS5jZnuSDkvz9wSFuxeDC25Z/S8RGha8rYrmK51EyEoxBrRiS+RcGh7JczLTi4aY
VMISaZavgWt3IprCX0ygJPdB1irSJHdeLsQ+lyBRNc3HLB3uQksSI5wzYZ++Fy+aGUEv9I07vWlg
zNyF0KMWvYogeRHWj2Edrvg1kDm7lKugizTbkIjggW8hyx81LSLWr1J2k3z5+epguPYSkp4PVUGn
hLJKwGBO0+ck0URXSf1fNj1JGEZENRlIxXuVuYajNmI85wbMtgb9hZUbw0QdiMyW1TteW05jgsZb
87BtzgbKcTtUuYaj4Yyb8OPyh86yLsVxnVh0YiHXMEWbpypSMraeS6SDnt3ReV8CyjXWnOaaXc0I
KlH6PPseSi73Zah2/AQ5vIcoBhsp+HbkFsCwOBhCFFfmOIezf3jJ2M7VYUZz4KQhePjgBz98gxDJ
a0gBo5xjPC2p1KYPgZVtsRfHNdUT27mSw52yMVzDa5EQfs6WHbfqeXYZW6lPQx5/+fnQu/EChxvA
dAr+XalEab7d0VNVGG5b4k5e1gAzF2ssKMBS33Sv4Ncw0pMl225LMCGrqwsAgEl/+dkALFGSbseY
XHfFx0C/+y/FrMAG8QQ3aZgTPLRGZohS7ad4dnCwy7i4OxYTmfLQyvcz3vPROOKIa0MWy/71qZsX
EvyW4D/r84MqMzUP80NHQMrXBsqh7HnOdtqpZGTrTsZeSBo3zRwVPxqoCu9F4YxDco75IONQYj1d
+yAEeu9DxOR+Q1B/yNW2VknzqgXRUMItuOnTaR7bghIiYIrF2AGL4EPnCiZ2XKtMTGTHAg1f1Baa
QSoKzIdmDkdgK1r/RwfvZzsYBw2BzzU++Seb8iPrBie0ff+tYZJyCNWMJKLlYWdDSsDm/YvHIX/e
9q2t8UyDSMchwR5qyrofYvIRFLPYO+69t/P0z6R+jLxPiJ9Wlqi+taNW6c+DqLb5hufl3IR4NcDd
QPV2WowiV9o40KMn6Q/mME1BfjDkVwD0bSzzlWLZfEaqWPSKGabMjlLs6KI59v5VimA7AMQnmBS5
H4z8XK+JbLxKOEzh8pc1k+iRV/ha3ggSrNO5ps0oyapkIuENlQQcjHJyMVxNbhNPgB+hwcP79bbr
XqvfHrc8n1wGDqJPG5L0tNROBAgHT5BHA2oIxnpYF2RDEasBC9KZFstss+JHpSHjPr7T3AAe72Vp
hN0pbWB2GmUDbhjHFUq3lYcHQS3odX6FfCzk+cl3mB8UhEMq6YD0shOFa4vk2gOxBgOEclcNjP12
5ENVPYPN5Hn0KitAhLy8s60T0zS7WFVVfIb8PhocM1HJ4pAKx9N86VFFZwO5y0AX+6OKacHtzp1W
tzqvJjF63k2cl+BFiaoxpTl6PgCO6OWL+HAQVsvpvxgJkBQpvQrnldwyYoimckcVX6GGAgpKSXyI
gFfrucdXm6mcHMA+rn/TtcM6/RALjx22UPiaiZmXCtuxmmXn2KT480Fmz4fKPRR58RDB2HeL5qi6
sYAdjZgtItWzga8RaMn6xZ0ANwdSbizznO8cTIz4Oreywdxlvl8j6NcSI35rTcPpSj70F2JNBK93
q7mQgAnoaqzUenSuIZkz7yQokckohE315RsRGSpR6d2xqLw8JiguFlLBQKChtHugoQG6pDkAFeGR
qON6+scWgMvhIww6OeasRH//xgk+I9JqOK6noaZCDyMxGThLZF8jl8wQ3RU3CLMfDGE48Tdk9dCD
Te55zwakePjjIF0d2qMRx9xQzyNkkxoGcJJTYy+RLulSstkHuPK6TzCufv5ZGcMs0CLZwK/iJVaL
xKPXaUByOffzCGxrXh+C6T9F5hd4AT2hxiMqX1xdVozE55Jtoc3ceIIyzwlxaHR1VpGFVWNKIrRo
1rmvMFUwNYKz6y+EP0x78JNedXwTWC+dSEaWcMNiHlqhPuvI8uVjgFyVnJocBHEUvhbSwxPlpSOl
ScTnGTIcNEOazB7NRFOz/kSKJ+ULXnDqAJy8ct57KesdTuWZefa1ofGccrdjy43gdwPE/+B4dxuI
IpKpfvZYS/KuGT7W74QO9cjiSHXOl4haITHCNQJ2v55nbaSexyv1Zu+OG3XCKlzlMtK1KnbnB+Kg
3SsvB78OaotZSydD5vGmjnV1KBLK0EEzdTP5I1aF1/dfdWifRcYSy/vwXrivciA0jGF97CCp1jAf
uVSal62rW2bkv186auuNTw9e0Kgr8UmHT7tahCmTFORxypaxF5Cp5dXM8cjeTPtPi4D1S+0kWHX/
ug7EoG78CvSj1mLWjIA/B62reDe4EGeeFNnNC2UyIKXDYthV+Eq3o0BQ3pKz9q0BNo5RGAPR6Vd5
EFRLz2GNRbx4yMryKk1mlhFIntkHP/BiiU/bvhydjyQgvcB8k2UP9zBTNhPdl2GjULAnB7XASdh5
dO4thGJJ0utRARMGT7UO8dWa1IP2hSQQ81gpORN+/5z7gqhwd6kpGM69fELPQ7l9NxKxowB4/XVG
zGaQw3MBg240BU1X+AHPVy/E+Le5OYPB9nhJSwfsEgTn3+kQn6BqlZ2pR7rNt3reWZltekzNRlae
qzuH31SIK3JyM/Uk/AODpS1KfDmYY8X2XHMOKuevmlDaEao1RERKOK6QoEh+fCynaDoNkWyaqi5g
3mvHmpPUmxlZDLD76xdcZPwiKyIPr2trL0kK+r3gQvtZrxH+M/+FsEYiUs0JHAR5V/Iq1SKMniiY
Ctg9TCYvK/CVwCfSEAtnF0P+j8ZiH1XmGC3M1d22JV+HnCQ+AmChQBerqOR+dehwo/8jEL7cljIt
Ah/3neH0zNZiXIXCB4rHsb5P2L4cfc6M8MbfUxwWAzTDOM8ifqtd8nj+eAOipGgVA3zY9V3mVCKr
3h8/9xZbZ8SZJQmRoAKZFjWoqJsi/0WYPUeWF1g31SrWLl8lpTz4rjrNgrSMAPbGfKYG0UcVs5Vf
q5GoQRHd+RNEjjhsi9NIgZrKB0nEg55U9dBgwIvRGEXLNPp8sC4qdErbBplpOODL6UX2E4K553hI
poCoE4ZDNRRvDaXDYiBSQvrtERLNXo98kw1FVelvizUJVNnCy8LwINV2MTti/6TBXd4X07Ya0GIV
8Mu3fny/J5E6hMxBeBjpyozrqzX5cVmDRncwo6V9OBT0gzI1qLnvv/z03sNB43csIurZK8+v0xoW
WVsNE/gHSc3rHXPZnr6MfY1vVrqS3/tSFKnUBc1uWBBaRkWFO1yIe1jsILqUEamB+Lq+Kcw71G8g
nmsP/RIMBesnxMrTbT94yYsnNiZ8ddSz6QVTtQbZsk3ijOaE64lQa8PZBMuVtN0I9CcJnWGcMMEe
c9s6wqqhY5uCIT9HtB2pwrgy6kZ8jpyu+Ge1NbiTTgAannHcyBVvGROMGNU0J8LGMr+MV8DA+6XG
RVxuC3DEaIEWKUvd08dm70HJMxKZk3eXDNlzRF+Zkh5WdUtlHK2qjmNd3UQ2XPO8vLLzIMt0BpzX
/Z4E6XoG4A58v3vR2b+a46og9cZiZbc5M/73nW/vC01pDWTfqlbHY1NHajFkcgz4GR56dyNIDNUv
KeAttz5cBMILqwstt3iBn8S1Zvi00zFyKsLx/AXpwkw9cuKyNQq5l/XrQcGZwU9q8lrK19Iunsvd
zzmkwpbBtVUjKI+ccO/yzRdn+P1yYASWvV8C1ISopgepadws8KaOYMi/dfDjLouFehYTZ3tJcBpP
RbcxmOeoo9QAbMHEddV/xUP7n8AqZAxNrh69iFLeA3ZnBJd6v3csv7frbHrEfVrnx+A9LJyMmhBx
OZ7Xz9U0r4TeDVHOxd9jFHp8F1BKONqjY5svCEyYJvi0fONvd1rO3gZc1kAPdqQcWEdJAYhErD+i
7ZlmMiaxRlhKXr/7Uc6EUZ1wItuAE7mz848rnjf5qfV3831096aZlsxi/jlN/1fxlQX17nX5RUyM
fpn4AwrYsNyrgk1zLIBusTjZzhYHFTwL1urbc9ncIRMrAE4d47wX4VLvEECf2MgJV8PESj0dEPL4
KfJMmhXuY32G+rhHmXV8QSRz6oIQdTs5A0bb3r2U8S29VhhV3I0vwQ/w5grS1juA5/Zg8e1Vzgkf
HzyNAG1F1efFzUdEwIzQ8pdnCJ5T1dWFBXn9Hk2gp0bVglX9W4XChfc5YQboscI5riBm2gUZa/mj
Z9kerEsRwQmePqTqi5b4m+r9y7DidG8eDPv2RUoOzjr5U0FG9rd+pZVhqLWuGyTrX1P2fcwZZGCW
mino11orUA6WXzxC7fynxMzGKieu9qMmYUYpIIwdjol4SPRzMimj2O0WsxA/RzX1eHYDzPW1nsrB
leihQ1jKZDryBfO+nZMYugF0VZBmuIMtWjMnInzsnqLTiVemWoMNj2rVQx2C3l0BxIAAe+Y0a+6G
QoLwbcsOm83A8jWbep82PR/bABFDLJcYGhzoXTT2YHfIIJZnwv8Jlgijx23UUjpsRWO/zFCYbENL
3QaxxjpqOLK1XszhxrlmUABhRM1TsntRGPzi6MBNQpRK0R9AvJ94ZCm7LqES3AID9g8prN4Qu1lt
JaxhBe8B39M63+vAlgluQbOw5Tb/WNpsT6WdoyQBtwwJXRn8F1ei2K7RhfvifOiM2nRhx9dI/Dx+
v97nwQXbFBc/CLfmASayiQDd9ohiy5GIKxihExoNinvlusdPGlWU4dPGl97AsgVbuFzgQ19eNLub
523QybXo6JVLdQzeKcoQeLlS61E/zEGX0BTOveNnY/nQLlOegFkWT/Wjy7tVpHNcZkIWH5H6evey
0o/8cSTIZP+NDFpZqt9GxREHpWLssMNaAYNxtx5SYWsRlkRJOJ9YGKJ7EsDFSEEUNDQ/Ly1Oxl9X
ZxizA3e+bMaag2PEwdu6Gzk4ymqf4ZhxKY4vLRkWBJMncDuqG8Ui1RqKBe/FKseYEHm+SwadPMav
Utwkwa43kMZMBNzQ+9m2Dv7wZcS/W50qDzNCyWNEBDzWMqO0gu7xtpHPqa3ihOQneDwfUnNiy7oS
mugH3bg3Fzdrj0BwyIxJqmXu/OO5vGtKRdzA637N+RWms86h0L7mjYx+eibBgFfeCQKcEg6iM6os
fWF10q0fPwKRnYn8yqO66fskA6u3EVQWJ+SvOpOP7UYHhrplDM3b0jnPUO2SKuvl5SGq4WFCwZq+
MpONtoIHi+mGbcWmL6TGf/4/mvNJRGQbLuFkzqqSIs45URRK//FWrs0YGJHz+fbdxEIEt+JgHnNx
kyvZsmRzmMMED6dZhgMzvcX9jW1i5u+iAKy1CbUGeLrPDtEnSzuBLLqJXA6kz3bBuZ1RVv9SpUU/
Lf+IZM0VhpkUbetOMt2HndWiOTugPm+py1hkX7w3yMfn9Keu/h5Dqa8JuAsEiX6I9WKgWvn9/lBU
bNwhrTTaEPctA+erzMj8w752i7L0TN85v6PMfADFNRsLMLnT47TcrHMas0ZNdP79OSFhDHEoNWf0
ugpmJvI1R53hG2TsMtlTR1xDjawyim+doRb5wJuSADNhSuBCHDCWms26jbUT9d/irkSpc2RzEQPt
7p33Yo+B0ckEVaZekWYV6XDxo+R7L6GIMpyc3dG8xLM7EdNxKe+JsCgeBt5Zq4sAsEmPBvBk/gDY
Lu6u2il7SQAmXz3dzXy9UgvVbs2EgBsVEn8PZEPjN+eMOHmDOVzZK9cKEcDt9AB1jd0nbkZ5gf73
yzboVXukcZqhjvAjKI3qYRAkIIxSkl99jlvYslhdNfq/iotzLAXXpXhN+xdJEXQhXqwnVKK3CCvs
lriXgOj7gXDUriwUDUCn4Sm67OBHyEESj1YuSQipi/sMY/4vRtrCH4ohlyBadsU2UB0oWxLxxl86
koUuCDPdorCp8xurN0kpHTYyOyLUEy0tCuT3UhPs+yn6Kz4jesbwfrCjPqQt1a59kaXwY52zwqR6
XHni9iat5OKsegIHSyAi/qG46WjDgFJHQKCIzpl86YGAqsE3UqR9+T32x1bw1azI52aKpvFkAV3G
uPnAcfe/RX3FPzAY7Mw5OTRsLst/rM/09ut8K6wdXZ/yOGOzLb6E+XLB511sH5V3Q+rGHAjnbBsz
9EcCwBx1BHX2F4KZMM3AoURxug+iWeo4Cw0DiolmWUYKL0mGqVKpbh/N80XCYjFIi2ZJPPIjqgKk
fTbIMXVddbJuoI5bhXjMaBeQoGZdLYEenBHwuO5Cww4CbPCH9WP6vt2cCPKG60o+lwHluPwu+P9c
C+7bGgGNSW5QocAEUBe5rD4FhtzpVBfPPonpf4K5JQgR3J5RIi78ZnmEhhQ6W48Ht9atywPt7tgJ
w6hIV900aCKYfa6PeCZg4yYWAB/KMuUUEPwYzaBsyHNyLAgQ3oBQFuE35ecjUBYHy2T91HRLdlzl
o/TiYWiBbu3Z1Y8dEOyF9zsqGNAAoGPzOkwhRJyVoAD2dkwWBAtu9HqF6XdS3YBY3reLjRXRCxdG
lmu67pKvJTTd9xyq0VwFcC5MRTzQ4w4n+E3hnWOkro2Su3gc3moXmznf6kAx3OwDRf/hzqvUZbCC
ArNSbmEQOIOkfIOOzkV2FAMzFmyKg0JK6r7FgXHgJABoZLzjw26Da4WSzC8is3AhK7PWgFiO4jT7
fe5Qj/I+bevXOMHeQIneMRL4YiJzr8o1FUvN7zPC+xN5hH/UzIMzlHOB9lH8773B/30y9Z2Optav
Gg3lJuqeN4R9X4uoryAst25FdKRe5YauwV9SL6jP8a9tzpPb0bUoJ13xvFCMgOCakMMi6+9PiRXM
t9Ym0Suv93QNsldMRJpt30kl2HCAmlzIgCXUKfOmBUGDVhCPVuZlUhRAUHlbvwLvBbur5FzEV8+3
3uDJ4WREO6AlqGI+1Ck7+FkCk23kgvDy3nd68GVM1/uoa9P7jPsFIqGx+F2a8BzweRlpOCVLQGI9
4d61LywyJC2ijaE+BAE9hRy1cQslCu6QoaYnUoTbFBbqiSQzPCEASlczyTA24OH1cbl79KYBSHSX
beS6l/a+URn+/FYuSONj51V3ZQ9jyYhT5rJ0YjKNpXZ7PQJKdp2CAiosxjKBt6kiDmNrHTj4UTwW
6sk9dlLM02nAr17AP7ASrKLfYOm+QrooPKhNT9xbIxoQeagc8acJ+WxrQNUDh7GRfa0XkfBKP1V2
ycIHRpiRgjV8DGbmvo8Y0dJ3hhiaxcjkaOgtI1XvkEr9CB3ZsemGS7PYXghAfXj3iigPSGATGPHL
/NxE8SkrmCO80TOVS1EhCnE6YTMfQMrK8o5+QZT11wo0RmkctWQRLMBTPGAG4bE6HHJzRZfWCwLV
FfOhtNhBuctva5vUOG6IL26azsxZj5SZbsU1POHuTu3E3pBRDrxcl0DfWHvIDUvWPY9PGAiCeHJu
k8ndJdZ3DXj69qKUISxyP6KYeBCoUBAngmN0G+2sYu/NHKX1effwlmsSGTDidNOPl54oqTeinR2Y
qJL2XXcAtFYHlFKuXELv2Kdz3wOjL7FHi5tqmuhw9VB5BxYUsLy8UmgNIoSuCIyoVSxbm4pE3m5x
qN8g3XQixyL2jJZ27xE0WQbxpHek+S8o3XDpbSvgtfLQlBtiUs9+xiWvZ0JBL7FwMmX7lqyJB8sO
eAoVqASHXQf5m1kggfCVgybIjy5K9L9BTd+YO7EZnfN70TslRsP9gYThEQI20uSZVh835Rc5I9C2
sKM5aLWWn4OkrQ8RD/vmeMnMoMNaW8y8p5r3jwBy+7Ff2ztz+Yk4LG7eEJUqyZiaIVKVMVlSNuoM
GUf6UYCxObg5reHsLgQyt1FEVGaIVou/2hH4ou45y6TqYpY21+trCMQSYPyVgjITocMnTJ6Wq3ik
Aumi1YZQEq871N1R4fDpIOkD3fWA4GH/jluDKUHFQ9xgIMk+jmhoXRWp0z2EV7nwnevu/r3Mh17i
9CCtVJd2AcxR+qNCjp9g6rrDsoiCJA7D+rG7YJsXG7c378Ve3gcLuRQ3mCRNvJim/p2BY1Yvxblk
TM2cf461ay2gAZr78uxTxPMIPbxLMfghDV89gQcxbEmz4CDE5jr4LcZwTXPHGrCagfpBDDJnj2Y4
Qqqq9Vtk1gP1ZQRjtgZKn6sK9cRmVJsIzaXC6iVHf1EFXC6VLqIZkdpVwrU6mCSaWcBAMMKWpgqt
BM1sgEPRgzmqagru98F5N1fcNSlPs9OFCce+kH6YoEBC2G7JZkvnjvEiSt1yw/mG7J0s22kYTRQc
sp657lLwNqopSDmFRtps0DjsuPVRfU1pSBXMWwtOgFIlbZ+MLyyx+Gi89ivKSbWl0B3nurYCHSuU
nIfjm8AyAybGIv4GgBjWNLAOQ8whV4M2ld7QHXB9PrRENct2YV8FmDmuCrMLkvczSc2zcbCfuajx
y5ia8WXVR7s5DwMhhX630q+8KRLUDX2Za+ZebvhXrPTyC0YSf6fZe3vYv9XbTMHqPbNybJXjQM04
KsJGcAjSHug3e/d2yhPRgbUa6m4fjuozo/RFisIv9fnVsmIKdBGIPMYrSS7SFNDAauqQB95rawfF
1ijxzBvmLCjcvcVzL/FDE6iKb6vJSXu0bvJs6dEgTy9/diW5fFjcfu4LsRNyJ4XGIF5ecj/wXnos
1NXHS0SmaKoQlDikvPQIlPP4zEVAK8om7F+kuGhURf2JDmPyC1DODwLQnxJZYo+Pz5R5kbspJ1A7
TlFeqvIoPPEx5hc9eDLBB6LjVbgQbDlCSmpILeVy2wxF0lgZ2vrJZbA0KXE8wJDZnKMH2xu6NFNN
BNRv8d2SmvZX5YrI8MKqsHT/7HXj8FflCZjGyJefsS1cx/XAVBNw9sQD0tAN+5pyCy8jASL6pig5
TXM5sNtUqNyw1PNp8eCHf16XFshGQG2DXqvbmni7P8ZqbawztKCX5qUjrs5JF42IMZabEpPpJ2NU
lkm2xYTndpMpVMd4Oy1g8Y05lyxNDpuaEetHzOrd1cEWY1SSJRElWWJUDjQveYfMoSUMogS9uh+9
bUkB92gdjFGL6obiSN/ccrkqQHJ5+NqlJviKeePwOskM3UavFHEg1E/4dfBS4th//XPOzPi4k9QH
hgXKCgGWrdS5S+WYGNP6k8RBDypOi+Voa/hwQsunzZdLe8RC/2mxtSSg4NRO8UdIvetwIbyLejJv
AjWt8CZoZ32oqKB6+lsid1ImkH/kJ6UJdB+07M9qsrWjMZ9ZeFzNw17QeyAiRFrXpOmmP/5o0ze4
khGUI0GFRP+ACcEruCsMe9Gd567vUU1+F6qw7GDeSUl2oa8d70gi/fnAKe97ONKQ2pP1L+DqYiwU
BDH3XZwESd7pZUEGg+DnCK8eg0q3hvOdl9Icw7ErjMFn8ytQldAKqOcC1pkMN0MEfSHHYn/pfXiz
EKVG3AErCrw/EHfqOwxx6WBn1ijkqFd1AoyZEYV17hG0ZUw5447z4j517yaCUNGFNgzwweR28g8j
KCSa5GLjB1mWIVsR/u1gbwOVUzw+OpxeLf9opoYZg9bZgZw8W6sL5cULnIt426o7vhpoQPHW2jRF
KZc6jYKt9bTaqzdY8fBH/Pf7aTdyClCHLdvDYmxf13IJfFWxY3qoYRkRSSWPG4v3X4moxRLAdetT
dVaUYnSEe5EkQyVmOpJ8QCGNXKcGr8Y/i4H69Kzk+rJKumiQbDsSDZliQPDM8vha3/5iGC/RC0cD
mi8reViNm0EjzWl8LTWH2Z6/OZbkpSV/15bi4xiOQp6Zk0iR8GUt46CbKpjVipdE27mQTN2pr8aq
owsftXvh+4rXkWYNmxRTVh4rN9HM3VKHHSrCkNlEPimE+Nl7Ne8mfTG6KYgkYjO4zUO6M1TKxBxf
dIFuA/uRJyCZBRLuG4ljl6lUeuUt3buUgATZKb4N5cgbFBfC4sGmPk+AxpYGp1+5V62TmJe3GYNt
7jJ1MqW82ICS3R5W8rWv/M2dEso1Mg7XXwBQWEmDokLQUEQiPULLgdrDeggWDgNexs3UnV67bbM2
VXF5wwyUMEif4Lmp69YZvg/tg+B7MU+mxvPBSMTg5GjOebUoQz7uJ+b7+FkZ3UNMigtMfg89omhB
hW4p+UZu7aVNrCwDzDHfwGdlKccAH4Ldd6iNKCcRL/GbR3a8PAABkncCikEQY8ijPP++Hhc9Ck9X
u5Xpndz1Cpdg0Bb1StJj/0+hYvL2mIyoDta7XOYR8Rei8dH2xMmSfqXQnR1+qDQ9vRHMq/scqoHx
zW4Tww5Uc4OR3pOH7DNfiBV5ba+wRGJO16f++l9bBQpujcdwTfJvQ7ouFZO6sdPb7zgVbxbiUa0U
sv+hevEECwrdeeEgopLQaK40U9MUTOujhykUka8L7+XoSKhikPCFRCmGF3EJJodMXxP+WTGggMnj
L2MDfNCp5amIhI11SgTfvOshfdigJDcDr3HrqZNIGgS4dJUcMwb06KD4jh+4Mjq4/UvLFo4/EZxy
GmATsptkTC3S2Xg8GuNI05wmNFoiQNZRu1CSL10lzj7P6aExkYmFUt2HBVCihmoOwixLF39xQqdr
uoAeKJwLHXB4I7DQkS5UcHBl48o7d6TK0pH1Pik3boIuD8quGQ11uqDKXU/kAy/ptIAK5LzS5off
vvFijDSFhm6Ladq0YihlCRh+MKfoiYTNU3o4DTOYds/O55CMz+Xquiitf4zioWxJj0tHrOF4k1wJ
2Li2OwnYW4JVoPz489ljl/XBJY7QLGm7qhx0G70FTjFDsSXwlFgRWQJIEvilMNXgeLvVcMzAA5XO
MVwble6NOPRMINOBE21lqXIYHnlK0D4qaOl0ZGGe5HPlceuuloZ6n5Y6oK4LeyStPuPocr6Vwvlp
CFRFujRpLhxA2XI3KrIOgDejO3LsBnaMqsZo7bRfSfBf4d4KVcCigYNbYh+e6ASU6H95V7W4mQwj
vnoF0U48ngNuKq24p+vx5Mc1b1XZGzNvFnXS8YgVDie5IJdCZuN6OmYX8fKt1hfTdLxgEsEx4ZfK
TbTRCElx3orG9tnk/oOfmoxYNBod4Eo1+jhUXhgZ2dFROZeOwLapz+trppDZXmT5NfKc1WPRC7qg
R/nIScn/ah9pvVl8VbM1KPGa6ojHoN9Fc3ibbzwkYts6zPmIkuiSEH5IIQcTqdFnduHiMounj7CX
ZmmEXr6zzt2o0eZwZ20NghCDnqJCxLgebjjbYA52Lvq97rhlm0kzeaiIEURCF+qst7pVF90mJlKv
KiuAw5Z4BcMprluKTgwOmijYZpTCiIo8C4dhxf3yTwL+aoyH6acTWSv8pUWvnZSUkJ5Dl1rrTYvo
7TlipwTPV8fAsXX7ur/aLSKSLcae/p9xVx8DfTO7FYv/ds5B+4L5sfCwJsPqfPQnOq6lu5wiwig4
4chFHOApqn/2PFrOAD8GnBxqSUPaIEuWYrCaod5t6zRvH4r1clxOyOLcSN0s8qEIbJoau/4hKKas
lE4uURTVKwNOlhXh/RWO7g1aqJxTYiwPbs02xVeDBZXjOzJd1cebLWTgFcZx73g2JzL4pmXUcTc+
6JUxFCVoSOmjXnMU9FXrkL0Km0dP6iiu25WCQrDe0fpF6e8SSHlLokFjPibPI5c0/UYPdDd8R4Mt
ar9EJlT+GcIMLpj2EMEUbVHijhvE5NRj0fC75KU+Geni04pmG173T/sDFxCy/hLs2MC7BI9C+Ip5
Su5rvAJSToMtdRt+2BlPyDgKCclM2ueJUhFOJCfC1TpVHJd4UeHti9jEirJcD8ZbOAlyIZmfxq5s
x8hLPedeAhuGc0l8i/rXzHNHW5W0AT1cXVJ9ssGRiWySR9dA1W0htId3VHMLiIOap72ZOIRR+nky
Gv2Ni30JaW71VGDHAeoTLyOuZytPaBA1Q5+O4tLBVw2bmu3Z5N4lOIIC9R4nOF0/xgAEk9SrwLtK
veybB+e2BIeP7V6AxAZ04mf86X+uCp01498zO85t6NJwYZ6fItCRujHVnpAseHh6dGl7wwxzbTvU
3zaEvs8uXRyx8CYSJKAKcpJFgQ6k1D2GxtfG1K995m4v5Q3ua5kzgREEa211r7/qqVEJ4nHLcoFK
5eaBWaY/s1K24KRXcJ6yAs10rX4/DStOAQeMS27PsCtPRVvDCgnjEfZB5qqjIzMZPO66HG6ZFhij
iXtdqKQu+rp/ibUzISEtxUuIE9YsH2JEZq0ooLmeA8TvqrB//DVxjxa6R3IV5cHZWSw99zq+Offq
TW5cWHlN0aECrvpmYCKqEvCuBqBCK5ZpyFvqBvTKBmeJIuQw8C2A8CFfvVfUdC6h8wMhGtDDDRkO
8LNNPmmotJYcIxc/EEWX/6z/GAZaZIgMWmBK1gZtZ+RXEE999hCvafHlmBEbZHa03ScnnVD3s7s8
RMBZlSf+XdE9NRqozeBahuF3iJUVmFYYtTyrdBK9orehZc1qrXlfc0dGLVHSesoeF2AeNfWGhO3W
tzHKwOl/DA19Sp5lrqPLa9zA/j1WZ3rgJavB9KAAHJ1AZfcDEBZQLvsO4Ve+HdETKxnW4aZt9hBr
3c1Axl4A84yiKgDe9/75NixPmvofjkWZSAB09R67fplOY0u64evCjIQZAaG67Xv2glHhEdQ06Rih
ww0XVkZdakQgvT35JzJJN2dOxQASMCQnAnRmjHT2LwN209XfOQVTiOnMvKrkVtCL1hfcX14GWqAY
UzE+OOcBKv04lzvlZJc+luj7xFZaVfFg8FJ/BFJ4aEQN2YfIPnQCiXGKNxDpPQA+4awJHl6uzAA1
elBErMsU7o0KEYUiSpqEonGtJvxG1UK+XCiHgKuWszaoeMDLV5EtluS3eeZujkPqLXED4utkh3M0
8gk6xr2fPy5VX/ryb47zIdZxScQ3BKsdhCwv7PLGyaYfs3pCbHsf2nxvjDnSfxUsXC25ahbiUZwK
B+58g1XNCh+I41gu5Av+Abjp/VhHMAn2qKN9O2bNjnZvAmP6SOxL0ngolYBSeqdfy3MCS7vkTHCk
NO49eWe1CamJ71hc28opFJDzKNkMWabGtYz/heZFEzr87cU/O3lD+j+NlckG8qWVppoL+0uhCSae
g8RzVu4ZTuzXprn7lIEK/+IhC70UYGlaZh0pfzQI0p3bfyxlozjhB8Fwce224fSXVDEAgJG5TyTY
LdQtu6qScXMao06nMsWvBy3gCGWs72M2WPA8dj2sxiSATMOoWbqQsxL2i0pbT3Mjb424dzzEYojJ
va/qFCX/XjYBkYN34cmU2XGiAn0jEAXLFp6yXhsneaHn8x7ZVnlqEPYXnX92cc9qqmih3sDGhaW5
es7EKatR5W0sxANyjjLWkyZ1Ka7hpMK09kpEvgvNYWk3m5xVJhtagyoWRPhcwxB7ThabtW6YsrrP
KjymogH+9MU2W45dyhii7ubibopBc19tYpqrBj81y3j9GYj1WptpaqVJ+0T2jl5wpCJGbNJjuJIk
zaR/0nWME79J8WpPIAKBzBzpnlY3qQoBbm1Z1rrYBINod0CLuv/viXb6gKB7hnsA1ttPRKtIfCah
Pmb+Vm/UVqJb+LM+uZvM8c3LQzb+SYsGsokTprhnrnkqFuPuKNkgOvrGY5ZIIUurlOkKc9tFJyIs
QqqlcfpgJAtJ0GQAuk8mm0ZC5QpFMb1Mza90+hF0gs7W++Fi4euHExekEBLfwBr+bmm6nsPXJH4/
tDgN/xmZ7+yh1pQKrOT/OgAeRXh71dJeqc8o1UaNUPDzovl/UiXt/YqxhTqhV6Dcl/Wje+YMQB5d
WXCe2mi9+oIKClJVUmsTWowUuG/t2aoMhjJZudFJ4G5jYyDlRIVZRce5KAJeqvF0P2QQHUHroazc
o+I01nAy8yBEbcRGfe7DC1qQSs0OLOr/5kwTe8lpPkMCuzUppyDsTm8VH1qEihoTrWqkRBKEQGvW
e6Iw2Bs579VJsVixOMNcTJetk6nDXMX5KmHloeHZXGHGvGYvyfKbELkun6W/JK0Pga0I2o0iJ19F
GureuxzRXB8mNk0xqtGNoi5uYIvnwz9vDZvtoX/VQuq8J9LKWJsxUgSHrhFwe9ozv74dMDOREOWV
VxYNxK1IkHAH7sFr2vY2HlNBNbgnH2vnlqidRfKGdF8Yq3JPgvAQXet2HMsm52QP7E43lgxjz5JH
I59DbbOMQC1dhswSnxRhrKFiQ57N5Chu+VUptnvVwMCX6gytjt1oAEpNEHxoe9M5j9X8sXIlgcCx
ag/ffyjh/1a+AgJB0gQlXVsfB0MJtgJsBEwS3yzKtjKPAgP37S9C9Rcvb605U1lslNk8aXvsoAA1
JWHCxAqb+ewmJOF+3lBPb3zWXLmXlCJWi33JisElYxi1k5mAWIb5Ea+7ZOtzHQYST9YkA4TPBLez
8py+M11+xvueJuFwsgVVMCBRDNI0nMfGZfTuTEXZoPshX058UgkSohlXAVbbb+9ufhMDNXho9AUI
xkJAfnqn1sidiJaGAK+RwkuIKQ4dzJVSnLa+qGgL3FOkeGKRXbqsNo1vBC7Imq2Yq5BhkbCz8UOk
kfti+wKWtw1AUPE5OjfxNKBPNUumhrqb7R3d8IJau4tYjfgft+Xz45v2ZqZbI78OXXZgAe9TuqYu
U3tku/FTZQCGnONwTbpqNWE+xpjGWUbQrOW+p9Vtze4mm4kOdXNAVkEv5ASEliep8Tf82vPc1SjV
Xw0X0eqVfe/N2ALnfEWvG48LFRASs0mY0ujPgRagqNz5YB/mV1qyJBmTtwtfGxh39p52nUX040t5
JBJwDElI44fTf1WPQU7r46XHv6plQDX17XaHljZe26kHtBf0+J/myvF7XWFi2A18fYsQGUNuVVIU
MWOlaY3CIqRW4SQ0VknMsWs3s8BLbrI7miAXFfmbIGyPZjuiq7cvTTkNBuwJbWI6Y+cURxexPuX7
TWFbOyB8xYlsgEBqXuaJp7cb4wEaYK+UfKiN34qaFQPSM8aCTqcTGZXZuLTz4/yB2kdyHemauKmJ
3Ke/2CNlfUIVuqwVbluFKqzB0gerTHAEWsXgHKV5o1RWdQhzM8g1iuf0Ghfb3q+/a+N8DU4mOhYR
ykQrtp1ZN4/3Limi6dALXa8rgMTzDNBdyax4Lp5WkFRd8Nl3jOONBIh1E5hjZl0Nk0wcNiU8DRMb
RHhGsrATTEp6kjQ9JYTHL7iaZyv9g8KV+BpILhfrvCVUwvXX3kptBQ==
`pragma protect end_protected

