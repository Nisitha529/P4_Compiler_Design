method Action _routing_add_entry(RoutingReqT key, RoutingRspT val);
